ROM_inst : ROM PORT MAP (
		address	 => address_sig,
		inclock	 => inclock_sig,
		q	 => q_sig
	);
