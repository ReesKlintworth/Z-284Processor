mux_1_inst : mux_1 PORT MAP (
		data0	 => data0_sig,
		data1	 => data1_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
