ROM_inst : ROM PORT MAP (
		address	 => address_sig,
		q	 => q_sig
	);
