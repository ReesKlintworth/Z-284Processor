ROM_2_inst : ROM_2 PORT MAP (
		address	 => address_sig,
		inclock	 => inclock_sig,
		q	 => q_sig
	);
