lpm_rom0_inst : lpm_rom0 PORT MAP (
		address	 => address_sig,
		q	 => q_sig
	);
