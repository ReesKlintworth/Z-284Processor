RAM_inst : RAM PORT MAP (
		address	 => address_sig,
		data	 => data_sig,
		inclock	 => inclock_sig,
		we	 => we_sig,
		q	 => q_sig
	);
